/**
 * GPR - Grouping Registers
 * @module_name gpr
 * @author Yongting Chen <yongting.chen@ucdconnect.ie>
 */
module gpr (
  
);
  
endmodule