module ctrl_testbench ();
   
endmodule